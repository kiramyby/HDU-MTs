module cpu(
    clk, rst_n, 
)